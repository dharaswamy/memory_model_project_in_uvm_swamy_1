`define MEM_DEPTH 4